// Copyright (C) 2017  Clifford Wolf <clifford@symbioticeda.com>
//
// Permission to use, copy, modify, and/or distribute this software for any
// purpose with or without fee is hereby granted, provided that the above
// copyright notice and this permission notice appear in all copies.
//
// THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
// WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
// MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
// ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
// WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
// ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
// OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.

`include "jg_define.sv"

module rvfi_testbench (
	input clock, reset
);

	`RVFI_WIRES

`ifdef YOSYS
	assume property (reset == $initstate);
`endif

	reg [7:0] cycle_reg = 0;
	wire [7:0] cycle = reset ? 0: cycle_reg;

	always @(posedge clock) begin
		cycle_reg <= reset ? 1 : cycle_reg + (cycle_reg != 255);
	end


	wire [6:0] insn_funct7 = rvfi_insn[31:25];
	wire [4:0] insn_rs2    = rvfi_insn[24:20];
	wire [4:0] insn_rs1    = rvfi_insn[19:15];
	wire [2:0] insn_funct3 = rvfi_insn[14:12];
	wire [4:0] insn_rd     = rvfi_insn[11: 7];
	wire [6:0] insn_opcode = rvfi_insn[ 6: 0];
	  

	`RISCV_FORMAL_CHECKER checker_inst (
		.clock  (clock),
		.reset  (cycle < `RISCV_FORMAL_RESET_CYCLES), //important to reduce proof time
`ifdef RISCV_FORMAL_TRIG_CYCLE
		.trig   (cycle == `RISCV_FORMAL_TRIG_CYCLE),
`endif
`ifdef RISCV_FORMAL_CHECK_CYCLE
		.check  (cycle == `RISCV_FORMAL_CHECK_CYCLE),
`endif
		`RVFI_CONN
	);

	rvfi_wrapper wrapper (
		.clock (clock),
		.reset (reset),
		`RVFI_CONN
	);
endmodule
